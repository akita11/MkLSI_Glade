*******************************************************************************
* CDL netlist
*
* Library : StdCell
* Top Cell Name: dff
* View Name: extracted
* Netlist created: 7.2.2017
*******************************************************************************

*.SCALE METER
*.GLOBAL Vdd Gnd

*******************************************************************************
* Library Name: StdCell
* Cell Name:    dff
* View Name:    extracted
*******************************************************************************

.SUBCKT dff CK Q D QB
*.PININFO CK:B Q:B D:B QB:B

MM6 n11 n7 Gnd Gnd nch w=6e-06 l=2e-06 as=2.4e-11 ps=1.4e-05 ad=4.8e-11 pd=2.2e-05 $X=8.8e-05 $Y=2.7e-05
MM9 n12 Q Gnd Gnd nch w=6e-06 l=2e-06 as=3e-11 ps=2.6e-05 ad=2.4e-11 pd=2.2e-05 $X=0.000124 $Y=2.7e-05
MM4 n10 n7 Gnd Gnd nch w=6e-06 l=2e-06 as=3e-11 ps=2.6e-05 ad=1.8e-11 pd=1.8e-05 $X=5.4e-05 $Y=2.7e-05
MM20 n16 Q Vdd Vdd pch w=1.8e-05 l=2e-06 as=5.4e-11 ps=3e-05 ad=9e-11 pd=3.8e-05 $X=0.000124 $Y=7.6e-05
MM7 n11 CK QB Gnd nch w=6e-06 l=2e-06 as=5.4e-11 ps=4.2e-05 ad=1.2e-11 pd=1.4e-05 $X=9.4e-05 $Y=2.7e-05
MM13 n6 CK n13 Vdd pch w=1.8e-05 l=2e-06 as=7.2e-11 ps=3.4e-05 ad=1.08e-10 pd=4.2e-05 $X=3.2e-05 $Y=7.6e-05
MM5 n7 n6 Gnd Gnd nch w=6e-06 l=2e-06 as=2.4e-11 ps=2.2e-05 ad=3e-11 pd=2.6e-05 $X=6.6e-05 $Y=2.7e-05
MM2 n9 n8 n6 Gnd nch w=6e-06 l=2e-06 as=4.2e-11 ps=3.4e-05 ad=1.8e-11 pd=1.8e-05 $X=3e-05 $Y=2.7e-05
MM21 Q QB Vdd Vdd pch w=1.8e-05 l=2e-06 as=1.8e-10 ps=3.8e-05 ad=1.44e-10 pd=3.4e-05 $X=0.000136 $Y=7.6e-05
MM15 n14 n7 Vdd Vdd pch w=1.8e-05 l=2e-06 as=5.4e-11 ps=3e-05 ad=9e-11 pd=3.8e-05 $X=5.4e-05 $Y=7.6e-05
MM14 n14 n8 n6 Vdd pch w=1.8e-05 l=2e-06 as=1.08e-10 ps=4.2e-05 ad=5.4e-11 pd=3e-05 $X=4.6e-05 $Y=7.6e-05
MM8 QB n8 n12 Gnd nch w=6e-06 l=2e-06 as=2.4e-11 ps=2.2e-05 ad=5.4e-11 pd=4.2e-05 $X=0.000114 $Y=2.7e-05
MM3 n6 CK n10 Gnd nch w=6e-06 l=2e-06 as=1.8e-11 ps=1.8e-05 ad=4.2e-11 pd=3.4e-05 $X=4.6e-05 $Y=2.7e-05
MM19 n16 CK QB Vdd pch w=1.8e-05 l=2e-06 as=1.8e-10 ps=5.8e-05 ad=5.4e-11 pd=3e-05 $X=0.000116 $Y=7.6e-05
MM18 QB n8 n15 Vdd pch w=1.8e-05 l=2e-06 as=3.6e-11 ps=2.6e-05 ad=1.8e-10 pd=5.8e-05 $X=9.4e-05 $Y=7.6e-05
MM17 n15 n7 Vdd Vdd pch w=1.8e-05 l=2e-06 as=7.2e-11 ps=3.4e-05 ad=3.6e-11 pd=2.6e-05 $X=8.8e-05 $Y=7.6e-05
MM16 n7 n6 Vdd Vdd pch w=1.8e-05 l=2e-06 as=1.8e-10 ps=3.8e-05 ad=1.44e-10 pd=3.4e-05 $X=6.6e-05 $Y=7.6e-05
MM12 n13 D Vdd Vdd pch w=1.8e-05 l=2e-06 as=9e-11 ps=3.8e-05 ad=7.2e-11 pd=3.4e-05 $X=2.2e-05 $Y=7.6e-05
MM11 n8 CK Vdd Vdd pch w=1.8e-05 l=2e-06 as=7.2e-11 ps=3.4e-05 ad=9e-11 pd=3.8e-05 $X=1e-05 $Y=7.6e-05
MM0 n8 CK Gnd Gnd nch w=6e-06 l=2e-06 as=6e-11 ps=2.6e-05 ad=4.8e-11 pd=2.2e-05 $X=1e-05 $Y=2.7e-05
MM1 n9 D Gnd Gnd nch w=6e-06 l=2e-06 as=1.8e-11 ps=1.8e-05 ad=3e-11 pd=2.6e-05 $X=2.2e-05 $Y=2.7e-05
MM10 Q QB Gnd Gnd nch w=6e-06 l=2e-06 as=2.4e-11 ps=2.2e-05 ad=3e-11 pd=2.6e-05 $X=0.000136 $Y=2.7e-05
.ENDS
